module Or8way (input wire [7:0] a, output wire b);
  assign b= |a;
endmodule
    
